library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_misc.all;
library altera;
use altera.altera_primitives_components.all;

entity counter_sync_test is
port (
    clk     : in std_logic;
    clearHC : in std_logic;
	 clearVC : in std_logic;
	 enableHC	:	in std_logic;
	 count_value_HC	:	out	std_logic_vector (11 downto 0);
	 count_value_VC	:	out	std_logic_vector (11 downto 0)
);
end counter_sync_test;


architecture basic of counter_sync_test is

component counter_12_bit is 
port(
	clk		: 	in		std_logic;
	zero		:	in		std_logic;
	enable	:	in		std_logic;
	count_value	:	out	std_logic_vector (11 downto 0)
);
end component;

signal	count_value_HC_tmp	:	std_logic_vector (11 downto 0);
signal	count_value_VC_tmp	:	std_logic_vector (11 downto 0);

begin

--- Replace this with your code ---
HC	:	counter_12_bit port map(
	clk		=>		clk,
	zero		=>		clearHC,
	enable	=>		enableHC,
	count_value	=>	count_value_HC_tmp
);

Hv	:	counter_12_bit port map(
	clk		=>		clk,
	zero		=>		clearVC,
	enable	=>		NOT count_value_HC_tmp(0) AND NOT count_value_HC_tmp(2) AND NOT count_value_HC_tmp(4) 
						AND NOT count_value_HC_tmp(5) AND NOT count_value_HC_tmp(6) AND NOT count_value_HC_tmp(7) 
						AND NOT count_value_HC_tmp(8) AND NOT count_value_HC_tmp(9) AND NOT count_value_HC_tmp(10) 
						AND NOT count_value_HC_tmp(11)
						AND count_value_HC_tmp(3) AND count_value_HC_tmp(1),
	count_value	=>	count_value_VC_tmp
);

count_value_HC <= count_value_HC_tmp;
count_value_VC <= count_value_VC_tmp;

end basic;